`define INN_MEM

`define SYSMAP_BASE_ADDR0  20'h01000
`define SYSMAP_FLG0        5'b01100

`define SYSMAP_BASE_ADDR1  20'h01001
`define SYSMAP_FLG1        5'b01100

`define SYSMAP_BASE_ADDR2  20'hfffff
`define SYSMAP_FLG2        5'b00000

`define SYSMAP_BASE_ADDR3  20'hfffff
`define SYSMAP_FLG3        5'b00000

`define SYSMAP_BASE_ADDR4  20'hfffff
`define SYSMAP_FLG4        5'b00000

`define SYSMAP_BASE_ADDR5  20'hfffff
`define SYSMAP_FLG5        5'b00000

`define SYSMAP_BASE_ADDR6  20'hfffff
`define SYSMAP_FLG6        5'b00000

`define SYSMAP_BASE_ADDR7  20'hfffff 
`define SYSMAP_FLG7        5'b00000

